module memory(
    input wire [7:0] mem_addr,             // Memory address
    inout wire [7:0] mem_data,             // Memory data
    input wire write_mem,                  // Write enable signal
    input wire clock                       // Clock signal
);
// Memory logic will be added here later
endmodule